LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
ENTITY fourto16decoder IS
PORT ( w: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
En : IN STD_LOGIC ;
s : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)) ;
END fourto16decoder;
ARCHITECTURE Behavior OF fourto16decoder IS
SIGNAL Enw : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
Enw <= EN&w;
WITH Enw SELECT
s <= "0000000000000001" WHEN "10000",
	  "0000000000000010" WHEN "10001",
	  "0000000000000100" WHEN "10010",
	  "0000000000001000" WHEN "10011",
	  "0000000000010000" WHEN "10100",
	  "0000000000100000" WHEN "10101",
	  "0000000001000000" WHEN "10110",
	  "0000000010000000" WHEN "10111",
	  "0000000100000000" WHEN "11000",
	  "0000001000000000" WHEN "11001",
	  "0000010000000000" WHEN "11010",
	  "0000100000000000" WHEN "11011",
	  "0001000000000000" WHEN "11100",
	  "0010000000000000" WHEN "11101",
	  "0100000000000000" WHEN "11110",
	  "1000000000000000" WHEN "11111",
	  "0000000000000000" WHEN OTHERS ;
END Behavior ;